`timescale 1ps / 1ps

module ow_rx_tb;

reg tb_din;
reg tb_clk;
wire ow_rst;


ow_rx rxi(
    .clk(tb_clk),
    .rst(ow_rst),
    .din(tb_din)
);

ow_rst rsti(
    .clk(tb_clk),
    .rst(1'b0),
    .din(tb_din),
    .ow_rst(ow_rst)
);

initial
begin
	tb_din = 0;
	tb_clk = 0;
end

always
begin
	#5000 tb_clk <= ~tb_clk;
end

initial
begin
	#1 tb_din <= 1'b1;
	#13880000 tb_din <= 1'b1;
	#4320000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#15679999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3080000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8360000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#15640000 tb_din <= 1'b0;
	#13839999 tb_din <= 1'b1;
	#23040000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#15040000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#15040000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#2638000000 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#4319999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#15679999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3080000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#22559999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#2243520000 tb_din <= 1'b0;
	#13839999 tb_din <= 1'b1;
	#4320000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#22559999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8040000 tb_din <= 1'b0;
	#2039999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15119999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#20160000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#20119999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8040000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#15120000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15119999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#20120000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2919999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#1495160000 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#4319999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#1760000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#15679999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#13880000 tb_din <= 1'b1;
	#22600000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8040000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15120000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15119999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8040000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#15120000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2040000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15119999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7159999 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#20120000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#20120000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#1818359999 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#4320000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1679999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#15680000 tb_din <= 1'b0;
	#1679999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#20919999 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#22880000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7159999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7159999 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#15039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2919999 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#15040000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#15039999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#15040000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7200000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#1813440000 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
	#4319999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8360000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#15679999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#13839999 tb_din <= 1'b1;
	#22720000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2119999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#15119999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15080000 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7159999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7119999 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#20120000 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2960000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7199999 tb_din <= 1'b1;
	#2920000 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#15079999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#2080000 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8000000 tb_din <= 1'b0;
	#2079999 tb_din <= 1'b1;
	#8039999 tb_din <= 1'b0;
	#7120000 tb_din <= 1'b1;
	#2959999 tb_din <= 1'b0;
	#2120000 tb_din <= 1'b1;
	#7999999 tb_din <= 1'b0;
	#7160000 tb_din <= 1'b1;
	#1908680000 tb_din <= 1'b0;
	#13839999 tb_din <= 1'b1;
	#4320000 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#20919999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15679999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#1759999 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8360000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8359999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3079999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#1680000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6999999 tb_din <= 1'b1;
	#3120000 tb_din <= 1'b0;
	#6959999 tb_din <= 1'b1;
	#15639999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#1719999 tb_din <= 1'b1;
	#8400000 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#8399999 tb_din <= 1'b0;
	#7000000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#6960000 tb_din <= 1'b1;
	#3119999 tb_din <= 1'b0;
	#1720000 tb_din <= 1'b1;
	#20919999 tb_din <= 1'b0;
	#13840000 tb_din <= 1'b1;
end
endmodule
